-- @file gs_initial_guess.vhd
-- @brief Q2.30 LUT for range [1.0, 2.0)
-- Guesses are in range [1.0, 0.5)

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity gs_initial_guess is
    port (
        address   : in std_logic_vector(7 downto 0);
        guess_out : out std_logic_vector(31 downto 0)
    );
end entity;

architecture behavioral of gs_initial_guess is
begin
    process(address)
    begin
        case address is
            when x"00" => guess_out <= x"40000000";
            when x"01" => guess_out <= x"3FC03FC0";
            when x"02" => guess_out <= x"3F80FE03";
            when x"03" => guess_out <= x"3F423954";
            when x"04" => guess_out <= x"3F03F03F";
            when x"05" => guess_out <= x"3EC62159";
            when x"06" => guess_out <= x"3E88CB3C";
            when x"07" => guess_out <= x"3E4BEC88";
            when x"08" => guess_out <= x"3E0F83E0";
            when x"09" => guess_out <= x"3DD38FF0";
            when x"0A" => guess_out <= x"3D980F66";
            when x"0B" => guess_out <= x"3D5D00F5";
            when x"0C" => guess_out <= x"3D226357";
            when x"0D" => guess_out <= x"3CE8354B";
            when x"0E" => guess_out <= x"3CAE7592";
            when x"0F" => guess_out <= x"3C7522F3";
            when x"10" => guess_out <= x"3C3C3C3C";
            when x"11" => guess_out <= x"3C03C03C";
            when x"12" => guess_out <= x"3BCBADC7";
            when x"13" => guess_out <= x"3B9403B9";
            when x"14" => guess_out <= x"3B5CC0ED";
            when x"15" => guess_out <= x"3B25E446";
            when x"16" => guess_out <= x"3AEF6CA9";
            when x"17" => guess_out <= x"3AB95900";
            when x"18" => guess_out <= x"3A83A83A";
            when x"19" => guess_out <= x"3A4E5947";
            when x"1A" => guess_out <= x"3A196B1E";
            when x"1B" => guess_out <= x"39E4DCB8";
            when x"1C" => guess_out <= x"39B0AD12";
            when x"1D" => guess_out <= x"397CDB2C";
            when x"1E" => guess_out <= x"3949660A";
            when x"1F" => guess_out <= x"39164CB5";
            when x"20" => guess_out <= x"38E38E38";
            when x"21" => guess_out <= x"38B129A2";
            when x"22" => guess_out <= x"387F1E03";
            when x"23" => guess_out <= x"384D6A72";
            when x"24" => guess_out <= x"381C0E07";
            when x"25" => guess_out <= x"37EB07DD";
            when x"26" => guess_out <= x"37BA5713";
            when x"27" => guess_out <= x"3789FACB";
            when x"28" => guess_out <= x"3759F229";
            when x"29" => guess_out <= x"372A3C56";
            when x"2A" => guess_out <= x"36FAD87B";
            when x"2B" => guess_out <= x"36CBC5C7";
            when x"2C" => guess_out <= x"369D0369";
            when x"2D" => guess_out <= x"366E9095";
            when x"2E" => guess_out <= x"36406C80";
            when x"2F" => guess_out <= x"36129663";
            when x"30" => guess_out <= x"35E50D79";
            when x"31" => guess_out <= x"35B7D0FF";
            when x"32" => guess_out <= x"358AE035";
            when x"33" => guess_out <= x"355E3A5F";
            when x"34" => guess_out <= x"3531DEC0";
            when x"35" => guess_out <= x"3505CCA2";
            when x"36" => guess_out <= x"34DA034D";
            when x"37" => guess_out <= x"34AE820E";
            when x"38" => guess_out <= x"34834834";
            when x"39" => guess_out <= x"3458550F";
            when x"3A" => guess_out <= x"342DA7F2";
            when x"3B" => guess_out <= x"34034034";
            when x"3C" => guess_out <= x"33D91D2A";
            when x"3D" => guess_out <= x"33AF3E2E";
            when x"3E" => guess_out <= x"3385A29D";
            when x"3F" => guess_out <= x"335C49D4";
            when x"40" => guess_out <= x"33333333";
            when x"41" => guess_out <= x"330A5E1B";
            when x"42" => guess_out <= x"32E1C9F0";
            when x"43" => guess_out <= x"32B97617";
            when x"44" => guess_out <= x"329161F9";
            when x"45" => guess_out <= x"32698CFF";
            when x"46" => guess_out <= x"3241F693";
            when x"47" => guess_out <= x"321A9E24";
            when x"48" => guess_out <= x"31F3831F";
            when x"49" => guess_out <= x"31CCA4F5";
            when x"4A" => guess_out <= x"31A6031A";
            when x"4B" => guess_out <= x"317F9D00";
            when x"4C" => guess_out <= x"3159721E";
            when x"4D" => guess_out <= x"313381EC";
            when x"4E" => guess_out <= x"310DCBE1";
            when x"4F" => guess_out <= x"30E84F79";
            when x"50" => guess_out <= x"30C30C30";
            when x"51" => guess_out <= x"309E0184";
            when x"52" => guess_out <= x"30792EF5";
            when x"53" => guess_out <= x"30549403";
            when x"54" => guess_out <= x"30303030";
            when x"55" => guess_out <= x"300C0300";
            when x"56" => guess_out <= x"2FE80BFA";
            when x"57" => guess_out <= x"2FC44AA2";
            when x"58" => guess_out <= x"2FA0BE82";
            when x"59" => guess_out <= x"2F7D6724";
            when x"5A" => guess_out <= x"2F5A4411";
            when x"5B" => guess_out <= x"2F3754D7";
            when x"5C" => guess_out <= x"2F149902";
            when x"5D" => guess_out <= x"2EF21023";
            when x"5E" => guess_out <= x"2ECFB9C8";
            when x"5F" => guess_out <= x"2EAD9584";
            when x"60" => guess_out <= x"2E8BA2E8";
            when x"61" => guess_out <= x"2E69E18A";
            when x"62" => guess_out <= x"2E4850FE";
            when x"63" => guess_out <= x"2E26F0DB";
            when x"64" => guess_out <= x"2E05C0B8";
            when x"65" => guess_out <= x"2DE4C02D";
            when x"66" => guess_out <= x"2DC3EED6";
            when x"67" => guess_out <= x"2DA34C4D";
            when x"68" => guess_out <= x"2D82D82D";
            when x"69" => guess_out <= x"2D629215";
            when x"6A" => guess_out <= x"2D4279A2";
            when x"6B" => guess_out <= x"2D228E75";
            when x"6C" => guess_out <= x"2D02D02D";
            when x"6D" => guess_out <= x"2CE33E6C";
            when x"6E" => guess_out <= x"2CC3D8D4";
            when x"6F" => guess_out <= x"2CA49F0A";
            when x"70" => guess_out <= x"2C8590B2";
            when x"71" => guess_out <= x"2C66AD71";
            when x"72" => guess_out <= x"2C47F4EE";
            when x"73" => guess_out <= x"2C2966D0";
            when x"74" => guess_out <= x"2C0B02C0";
            when x"75" => guess_out <= x"2BECC868";
            when x"76" => guess_out <= x"2BCEB771";
            when x"77" => guess_out <= x"2BB0CF87";
            when x"78" => guess_out <= x"2B931057";
            when x"79" => guess_out <= x"2B75798C";
            when x"7A" => guess_out <= x"2B580AD6";
            when x"7B" => guess_out <= x"2B3AC3E2";
            when x"7C" => guess_out <= x"2B1DA461";
            when x"7D" => guess_out <= x"2B00AC02";
            when x"7E" => guess_out <= x"2AE3DA78";
            when x"7F" => guess_out <= x"2AC72F74";
            when x"80" => guess_out <= x"2AAAAAAA";
            when x"81" => guess_out <= x"2A8E4BCD";
            when x"82" => guess_out <= x"2A721291";
            when x"83" => guess_out <= x"2A55FEAD";
            when x"84" => guess_out <= x"2A3A0FD5";
            when x"85" => guess_out <= x"2A1E45C2";
            when x"86" => guess_out <= x"2A02A02A";
            when x"87" => guess_out <= x"29E71EC5";
            when x"88" => guess_out <= x"29CBC14E";
            when x"89" => guess_out <= x"29B0877D";
            when x"8A" => guess_out <= x"2995710E";
            when x"8B" => guess_out <= x"297A7DBB";
            when x"8C" => guess_out <= x"295FAD40";
            when x"8D" => guess_out <= x"2944FF5A";
            when x"8E" => guess_out <= x"292A73C7";
            when x"8F" => guess_out <= x"29100A44";
            when x"90" => guess_out <= x"28F5C28F";
            when x"91" => guess_out <= x"28DB9C68";
            when x"92" => guess_out <= x"28C1978F";
            when x"93" => guess_out <= x"28A7B3C5";
            when x"94" => guess_out <= x"288DF0CA";
            when x"95" => guess_out <= x"28744E61";
            when x"96" => guess_out <= x"285ACC4B";
            when x"97" => guess_out <= x"28416A4C";
            when x"98" => guess_out <= x"28282828";
            when x"99" => guess_out <= x"280F05A2";
            when x"9A" => guess_out <= x"27F6027F";
            when x"9B" => guess_out <= x"27DD1E85";
            when x"9C" => guess_out <= x"27C45979";
            when x"9D" => guess_out <= x"27ABB323";
            when x"9E" => guess_out <= x"27932B48";
            when x"9F" => guess_out <= x"277AC1B2";
            when x"A0" => guess_out <= x"27627627";
            when x"A1" => guess_out <= x"274A4870";
            when x"A2" => guess_out <= x"27323858";
            when x"A3" => guess_out <= x"271A45A6";
            when x"A4" => guess_out <= x"27027027";
            when x"A5" => guess_out <= x"26EAB7A3";
            when x"A6" => guess_out <= x"26D31BE7";
            when x"A7" => guess_out <= x"26BB9CBF";
            when x"A8" => guess_out <= x"26A439F6";
            when x"A9" => guess_out <= x"268CF359";
            when x"AA" => guess_out <= x"2675C8B6";
            when x"AB" => guess_out <= x"265EB9DA";
            when x"AC" => guess_out <= x"2647C694";
            when x"AD" => guess_out <= x"2630EEB1";
            when x"AE" => guess_out <= x"261A3202";
            when x"AF" => guess_out <= x"26039055";
            when x"B0" => guess_out <= x"25ED097B";
            when x"B1" => guess_out <= x"25D69D43";
            when x"B2" => guess_out <= x"25C04B80";
            when x"B3" => guess_out <= x"25AA1402";
            when x"B4" => guess_out <= x"2593F69B";
            when x"B5" => guess_out <= x"257DF31C";
            when x"B6" => guess_out <= x"2568095A";
            when x"B7" => guess_out <= x"25523925";
            when x"B8" => guess_out <= x"253C8253";
            when x"B9" => guess_out <= x"2526E4B7";
            when x"BA" => guess_out <= x"25116025";
            when x"BB" => guess_out <= x"24FBF471";
            when x"BC" => guess_out <= x"24E6A171";
            when x"BD" => guess_out <= x"24D166F9";
            when x"BE" => guess_out <= x"24BC44E1";
            when x"BF" => guess_out <= x"24A73AFD";
            when x"C0" => guess_out <= x"24924924";
            when x"C1" => guess_out <= x"247D6F2E";
            when x"C2" => guess_out <= x"2468ACF1";
            when x"C3" => guess_out <= x"24540245";
            when x"C4" => guess_out <= x"243F6F02";
            when x"C5" => guess_out <= x"242AF300";
            when x"C6" => guess_out <= x"24168E18";
            when x"C7" => guess_out <= x"24024024";
            when x"C8" => guess_out <= x"23EE08FB";
            when x"C9" => guess_out <= x"23D9E878";
            when x"CA" => guess_out <= x"23C5DE76";
            when x"CB" => guess_out <= x"23B1EACE";
            when x"CC" => guess_out <= x"239E0D5B";
            when x"CD" => guess_out <= x"238A45F8";
            when x"CE" => guess_out <= x"23769480";
            when x"CF" => guess_out <= x"2362F8CF";
            when x"D0" => guess_out <= x"234F72C2";
            when x"D1" => guess_out <= x"233C0233";
            when x"D2" => guess_out <= x"2328A701";
            when x"D3" => guess_out <= x"23156107";
            when x"D4" => guess_out <= x"23023023";
            when x"D5" => guess_out <= x"22EF1432";
            when x"D6" => guess_out <= x"22DC0D12";
            when x"D7" => guess_out <= x"22C91AA1";
            when x"D8" => guess_out <= x"22B63CBE";
            when x"D9" => guess_out <= x"22A37347";
            when x"DA" => guess_out <= x"2290BE1C";
            when x"DB" => guess_out <= x"227E1D1A";
            when x"DC" => guess_out <= x"226B9022";
            when x"DD" => guess_out <= x"22591713";
            when x"DE" => guess_out <= x"2246B1CE";
            when x"DF" => guess_out <= x"22346033";
            when x"E0" => guess_out <= x"22222222";
            when x"E1" => guess_out <= x"220FF77C";
            when x"E2" => guess_out <= x"21FDE021";
            when x"E3" => guess_out <= x"21EBDBF5";
            when x"E4" => guess_out <= x"21D9EAD7";
            when x"E5" => guess_out <= x"21C80CAB";
            when x"E6" => guess_out <= x"21B64151";
            when x"E7" => guess_out <= x"21A488AC";
            when x"E8" => guess_out <= x"2192E29F";
            when x"E9" => guess_out <= x"21814F0D";
            when x"EA" => guess_out <= x"216FCDD8";
            when x"EB" => guess_out <= x"215E5EE4";
            when x"EC" => guess_out <= x"214D0214";
            when x"ED" => guess_out <= x"213BB74D";
            when x"EE" => guess_out <= x"212A7E72";
            when x"EF" => guess_out <= x"21195766";
            when x"F0" => guess_out <= x"21084210";
            when x"F1" => guess_out <= x"20F73E53";
            when x"F2" => guess_out <= x"20E64C14";
            when x"F3" => guess_out <= x"20D56B38";
            when x"F4" => guess_out <= x"20C49BA5";
            when x"F5" => guess_out <= x"20B3DD40";
            when x"F6" => guess_out <= x"20A32FEF";
            when x"F7" => guess_out <= x"20929398";
            when x"F8" => guess_out <= x"20820820";
            when x"F9" => guess_out <= x"20718D6F";
            when x"FA" => guess_out <= x"2061236A";
            when x"FB" => guess_out <= x"2050C9F8";
            when x"FC" => guess_out <= x"20408102";
            when x"FD" => guess_out <= x"2030486C";
            when x"FE" => guess_out <= x"20202020";
            when x"FF" => guess_out <= x"20100804";
            when others => guess_out <= x"40000000";
        end case;
    end process;
end architecture;