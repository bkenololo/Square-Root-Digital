-- @file nr_initial_guess.vhd
-- @brief Q2.30 LUT for Sqrt(x) where x in [1.0, 2.0)
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity nr_initial_guess is
    port (address : in std_logic_vector(9 downto 0); initial_guess_out : out std_logic_vector(31 downto 0));
end entity;

architecture rtl of nr_initial_guess is
    type rom_type is array (0 to 1023) of std_logic_vector(31 downto 0);
    constant INITIAL_GUESS_TABLE : rom_type := (
        0 => x"40000000",
        1 => x"4007FF80",
        2 => x"400FFE00",
        3 => x"4017FB81",
        4 => x"401FF803",
        5 => x"4027F387",
        6 => x"402FEE0D",
        7 => x"4037E795",
        8 => x"403FE01F",
        9 => x"4047D7AD",
        10 => x"404FCE3E",
        11 => x"4057C3D2",
        12 => x"405FB86B",
        13 => x"4067AC08",
        14 => x"406F9EAA",
        15 => x"40779051",
        16 => x"407F80FD",
        17 => x"408770AF",
        18 => x"408F5F68",
        19 => x"40974D27",
        20 => x"409F39ED",
        21 => x"40A725BB",
        22 => x"40AF1090",
        23 => x"40B6FA6D",
        24 => x"40BEE353",
        25 => x"40C6CB41",
        26 => x"40CEB239",
        27 => x"40D6983A",
        28 => x"40DE7D44",
        29 => x"40E66159",
        30 => x"40EE4479",
        31 => x"40F626A3",
        32 => x"40FE07D8",
        33 => x"4105E819",
        34 => x"410DC766",
        35 => x"4115A5BF",
        36 => x"411D8325",
        37 => x"41255F98",
        38 => x"412D3B17",
        39 => x"413515A5",
        40 => x"413CEF40",
        41 => x"4144C7EA",
        42 => x"414C9FA3",
        43 => x"4154766A",
        44 => x"415C4C41",
        45 => x"41642127",
        46 => x"416BF51D",
        47 => x"4173C824",
        48 => x"417B9A3B",
        49 => x"41836B64",
        50 => x"418B3B9D",
        51 => x"41930AE9",
        52 => x"419AD946",
        53 => x"41A2A6B6",
        54 => x"41AA7338",
        55 => x"41B23ECD",
        56 => x"41BA0976",
        57 => x"41C1D332",
        58 => x"41C99C03",
        59 => x"41D163E7",
        60 => x"41D92AE1",
        61 => x"41E0F0EF",
        62 => x"41E8B612",
        63 => x"41F07A4B",
        64 => x"41F83D9A",
        65 => x"42000000",
        66 => x"4207C17B",
        67 => x"420F820E",
        68 => x"421741B8",
        69 => x"421F0079",
        70 => x"4226BE53",
        71 => x"422E7B44",
        72 => x"4236374E",
        73 => x"423DF271",
        74 => x"4245ACAD",
        75 => x"424D6602",
        76 => x"42551E71",
        77 => x"425CD5FB",
        78 => x"42648C9E",
        79 => x"426C425C",
        80 => x"4273F736",
        81 => x"427BAB2A",
        82 => x"42835E3B",
        83 => x"428B1067",
        84 => x"4292C1AF",
        85 => x"429A7214",
        86 => x"42A22196",
        87 => x"42A9D035",
        88 => x"42B17DF1",
        89 => x"42B92ACB",
        90 => x"42C0D6C4",
        91 => x"42C881DA",
        92 => x"42D02C10",
        93 => x"42D7D564",
        94 => x"42DF7DD8",
        95 => x"42E7256B",
        96 => x"42EECC1E",
        97 => x"42F671F2",
        98 => x"42FE16E5",
        99 => x"4305BAFA",
        100 => x"430D5E30",
        101 => x"43150087",
        102 => x"431CA200",
        103 => x"4324429B",
        104 => x"432BE258",
        105 => x"43338137",
        106 => x"433B1F3A",
        107 => x"4342BC60",
        108 => x"434A58A9",
        109 => x"4351F416",
        110 => x"43598EA7",
        111 => x"4361285C",
        112 => x"4368C136",
        113 => x"43705935",
        114 => x"4377F059",
        115 => x"437F86A2",
        116 => x"43871C11",
        117 => x"438EB0A7",
        118 => x"43964462",
        119 => x"439DD745",
        120 => x"43A5694E",
        121 => x"43ACFA7E",
        122 => x"43B48AD6",
        123 => x"43BC1A56",
        124 => x"43C3A8FE",
        125 => x"43CB36CE",
        126 => x"43D2C3C7",
        127 => x"43DA4FE8",
        128 => x"43E1DB33",
        129 => x"43E965A7",
        130 => x"43F0EF45",
        131 => x"43F8780D",
        132 => x"44000000",
        133 => x"4407871C",
        134 => x"440F0D64",
        135 => x"441692D7",
        136 => x"441E1775",
        137 => x"44259B3F",
        138 => x"442D1E35",
        139 => x"4434A057",
        140 => x"443C21A6",
        141 => x"4443A221",
        142 => x"444B21C9",
        143 => x"4452A09F",
        144 => x"445A1EA2",
        145 => x"44619BD3",
        146 => x"44691833",
        147 => x"447093C0",
        148 => x"44780E7D",
        149 => x"447F8868",
        150 => x"44870182",
        151 => x"448E79CC",
        152 => x"4495F146",
        153 => x"449D67EF",
        154 => x"44A4DDC9",
        155 => x"44AC52D3",
        156 => x"44B3C70F",
        157 => x"44BB3A7B",
        158 => x"44C2AD18",
        159 => x"44CA1EE7",
        160 => x"44D18FE8",
        161 => x"44D9001B",
        162 => x"44E06F81",
        163 => x"44E7DE19",
        164 => x"44EF4BE4",
        165 => x"44F6B8E2",
        166 => x"44FE2513",
        167 => x"45059078",
        168 => x"450CFB11",
        169 => x"451464DE",
        170 => x"451BCDE0",
        171 => x"45233616",
        172 => x"452A9D81",
        173 => x"45320422",
        174 => x"453969F7",
        175 => x"4540CF03",
        176 => x"45483344",
        177 => x"454F96BC",
        178 => x"4556F96A",
        179 => x"455E5B4F",
        180 => x"4565BC6B",
        181 => x"456D1CBE",
        182 => x"45747C48",
        183 => x"457BDB0A",
        184 => x"45833904",
        185 => x"458A9637",
        186 => x"4591F2A1",
        187 => x"45994E45",
        188 => x"45A0A921",
        189 => x"45A80337",
        190 => x"45AF5C86",
        191 => x"45B6B50E",
        192 => x"45BE0CD1",
        193 => x"45C563CE",
        194 => x"45CCBA05",
        195 => x"45D40F77",
        196 => x"45DB6424",
        197 => x"45E2B80C",
        198 => x"45EA0B2F",
        199 => x"45F15D8E",
        200 => x"45F8AF29",
        201 => x"46000000",
        202 => x"46075013",
        203 => x"460E9F63",
        204 => x"4615EDEF",
        205 => x"461D3BB9",
        206 => x"462488C0",
        207 => x"462BD505",
        208 => x"46332087",
        209 => x"463A6B47",
        210 => x"4641B546",
        211 => x"4648FE83",
        212 => x"465046FF",
        213 => x"46578EB9",
        214 => x"465ED5B3",
        215 => x"46661BED",
        216 => x"466D6166",
        217 => x"4674A61F",
        218 => x"467BEA18",
        219 => x"46832D51",
        220 => x"468A6FCB",
        221 => x"4691B186",
        222 => x"4698F282",
        223 => x"46A032BF",
        224 => x"46A7723D",
        225 => x"46AEB0FE",
        226 => x"46B5EF00",
        227 => x"46BD2C44",
        228 => x"46C468CB",
        229 => x"46CBA495",
        230 => x"46D2DFA1",
        231 => x"46DA19F1",
        232 => x"46E15383",
        233 => x"46E88C5A",
        234 => x"46EFC474",
        235 => x"46F6FBD2",
        236 => x"46FE3274",
        237 => x"4705685B",
        238 => x"470C9D86",
        239 => x"4713D1F7",
        240 => x"471B05AC",
        241 => x"472238A7",
        242 => x"47296AE7",
        243 => x"47309C6D",
        244 => x"4737CD3A",
        245 => x"473EFD4C",
        246 => x"47462CA5",
        247 => x"474D5B44",
        248 => x"4754892A",
        249 => x"475BB658",
        250 => x"4762E2CC",
        251 => x"476A0E88",
        252 => x"4771398C",
        253 => x"477863D8",
        254 => x"477F8D6C",
        255 => x"4786B649",
        256 => x"478DDE6E",
        257 => x"479505DC",
        258 => x"479C2C93",
        259 => x"47A35293",
        260 => x"47AA77DD",
        261 => x"47B19C70",
        262 => x"47B8C04D",
        263 => x"47BFE374",
        264 => x"47C705E6",
        265 => x"47CE27A2",
        266 => x"47D548A9",
        267 => x"47DC68FB",
        268 => x"47E38898",
        269 => x"47EAA780",
        270 => x"47F1C5B4",
        271 => x"47F8E334",
        272 => x"48000000",
        273 => x"48071C17",
        274 => x"480E377C",
        275 => x"4815522D",
        276 => x"481C6C2A",
        277 => x"48238575",
        278 => x"482A9E0D",
        279 => x"4831B5F3",
        280 => x"4838CD26",
        281 => x"483FE3A7",
        282 => x"4846F976",
        283 => x"484E0E93",
        284 => x"485522FF",
        285 => x"485C36B9",
        286 => x"486349C3",
        287 => x"486A5C1B",
        288 => x"48716DC3",
        289 => x"48787EBA",
        290 => x"487F8F01",
        291 => x"48869E98",
        292 => x"488DAD7E",
        293 => x"4894BBB6",
        294 => x"489BC93D",
        295 => x"48A2D615",
        296 => x"48A9E23F",
        297 => x"48B0EDB9",
        298 => x"48B7F884",
        299 => x"48BF02A1",
        300 => x"48C60C10",
        301 => x"48CD14D1",
        302 => x"48D41CE3",
        303 => x"48DB2448",
        304 => x"48E22B00",
        305 => x"48E9310A",
        306 => x"48F03667",
        307 => x"48F73B16",
        308 => x"48FE3F1A",
        309 => x"49054270",
        310 => x"490C451B",
        311 => x"49134719",
        312 => x"491A486B",
        313 => x"49214911",
        314 => x"4928490C",
        315 => x"492F485B",
        316 => x"493646FF",
        317 => x"493D44F9",
        318 => x"49444247",
        319 => x"494B3EEB",
        320 => x"49523AE4",
        321 => x"49593633",
        322 => x"496030D8",
        323 => x"49672AD3",
        324 => x"496E2424",
        325 => x"49751CCC",
        326 => x"497C14CB",
        327 => x"49830C20",
        328 => x"498A02CD",
        329 => x"4990F8D0",
        330 => x"4997EE2C",
        331 => x"499EE2DE",
        332 => x"49A5D6E9",
        333 => x"49ACCA4C",
        334 => x"49B3BD07",
        335 => x"49BAAF1A",
        336 => x"49C1A086",
        337 => x"49C8914A",
        338 => x"49CF8168",
        339 => x"49D670DE",
        340 => x"49DD5FAE",
        341 => x"49E44DD8",
        342 => x"49EB3B5B",
        343 => x"49F22837",
        344 => x"49F9146E",
        345 => x"4A000000",
        346 => x"4A06EAEB",
        347 => x"4A0DD531",
        348 => x"4A14BED2",
        349 => x"4A1BA7CE",
        350 => x"4A229025",
        351 => x"4A2977D7",
        352 => x"4A305EE4",
        353 => x"4A37454E",
        354 => x"4A3E2B13",
        355 => x"4A451034",
        356 => x"4A4BF4B1",
        357 => x"4A52D88B",
        358 => x"4A59BBC1",
        359 => x"4A609E54",
        360 => x"4A678044",
        361 => x"4A6E6191",
        362 => x"4A75423B",
        363 => x"4A7C2243",
        364 => x"4A8301A8",
        365 => x"4A89E06B",
        366 => x"4A90BE8C",
        367 => x"4A979C0B",
        368 => x"4A9E78E8",
        369 => x"4AA55524",
        370 => x"4AAC30BF",
        371 => x"4AB30BB8",
        372 => x"4AB9E610",
        373 => x"4AC0BFC8",
        374 => x"4AC798DF",
        375 => x"4ACE7155",
        376 => x"4AD5492B",
        377 => x"4ADC2061",
        378 => x"4AE2F6F7",
        379 => x"4AE9CCED",
        380 => x"4AF0A244",
        381 => x"4AF776FB",
        382 => x"4AFE4B12",
        383 => x"4B051E8B",
        384 => x"4B0BF165",
        385 => x"4B12C3A0",
        386 => x"4B19953C",
        387 => x"4B20663A",
        388 => x"4B27369A",
        389 => x"4B2E065B",
        390 => x"4B34D57F",
        391 => x"4B3BA405",
        392 => x"4B4271ED",
        393 => x"4B493F38",
        394 => x"4B500BE5",
        395 => x"4B56D7F6",
        396 => x"4B5DA369",
        397 => x"4B646E40",
        398 => x"4B6B387A",
        399 => x"4B720218",
        400 => x"4B78CB19",
        401 => x"4B7F937E",
        402 => x"4B865B48",
        403 => x"4B8D2275",
        404 => x"4B93E907",
        405 => x"4B9AAEFE",
        406 => x"4BA17459",
        407 => x"4BA83919",
        408 => x"4BAEFD3E",
        409 => x"4BB5C0C9",
        410 => x"4BBC83B8",
        411 => x"4BC3460D",
        412 => x"4BCA07C8",
        413 => x"4BD0C8E9",
        414 => x"4BD78970",
        415 => x"4BDE495D",
        416 => x"4BE508B0",
        417 => x"4BEBC76A",
        418 => x"4BF2858A",
        419 => x"4BF94311",
        420 => x"4C000000",
        421 => x"4C06BC55",
        422 => x"4C0D7811",
        423 => x"4C143335",
        424 => x"4C1AEDC1",
        425 => x"4C21A7B4",
        426 => x"4C286110",
        427 => x"4C2F19D3",
        428 => x"4C35D1FE",
        429 => x"4C3C8992",
        430 => x"4C43408F",
        431 => x"4C49F6F4",
        432 => x"4C50ACC2",
        433 => x"4C5761F9",
        434 => x"4C5E1699",
        435 => x"4C64CAA3",
        436 => x"4C6B7E16",
        437 => x"4C7230F3",
        438 => x"4C78E339",
        439 => x"4C7F94E9",
        440 => x"4C864604",
        441 => x"4C8CF689",
        442 => x"4C93A678",
        443 => x"4C9A55D1",
        444 => x"4CA10496",
        445 => x"4CA7B2C5",
        446 => x"4CAE605F",
        447 => x"4CB50D65",
        448 => x"4CBBB9D5",
        449 => x"4CC265B2",
        450 => x"4CC910F9",
        451 => x"4CCFBBAD",
        452 => x"4CD665CC",
        453 => x"4CDD0F58",
        454 => x"4CE3B850",
        455 => x"4CEA60B4",
        456 => x"4CF10884",
        457 => x"4CF7AFC2",
        458 => x"4CFE566C",
        459 => x"4D04FC83",
        460 => x"4D0BA207",
        461 => x"4D1246F9",
        462 => x"4D18EB58",
        463 => x"4D1F8F24",
        464 => x"4D26325E",
        465 => x"4D2CD506",
        466 => x"4D33771C",
        467 => x"4D3A18A0",
        468 => x"4D40B993",
        469 => x"4D4759F4",
        470 => x"4D4DF9C3",
        471 => x"4D549902",
        472 => x"4D5B37AF",
        473 => x"4D61D5CB",
        474 => x"4D687356",
        475 => x"4D6F1051",
        476 => x"4D75ACBB",
        477 => x"4D7C4894",
        478 => x"4D82E3DE",
        479 => x"4D897E97",
        480 => x"4D9018C1",
        481 => x"4D96B25A",
        482 => x"4D9D4B64",
        483 => x"4DA3E3DE",
        484 => x"4DAA7BC9",
        485 => x"4DB11325",
        486 => x"4DB7A9F2",
        487 => x"4DBE402F",
        488 => x"4DC4D5DE",
        489 => x"4DCB6AFE",
        490 => x"4DD1FF90",
        491 => x"4DD89393",
        492 => x"4DDF2708",
        493 => x"4DE5B9EF",
        494 => x"4DEC4C47",
        495 => x"4DF2DE12",
        496 => x"4DF96F50",
        497 => x"4E000000",
        498 => x"4E069022",
        499 => x"4E0D1FB7",
        500 => x"4E13AEBF",
        501 => x"4E1A3D3A",
        502 => x"4E20CB28",
        503 => x"4E275889",
        504 => x"4E2DE55E",
        505 => x"4E3471A6",
        506 => x"4E3AFD62",
        507 => x"4E418892",
        508 => x"4E481336",
        509 => x"4E4E9D4E",
        510 => x"4E5526DA",
        511 => x"4E5BAFDB",
        512 => x"4E623850",
        513 => x"4E68C039",
        514 => x"4E6F4798",
        515 => x"4E75CE6B",
        516 => x"4E7C54B4",
        517 => x"4E82DA71",
        518 => x"4E895FA4",
        519 => x"4E8FE44D",
        520 => x"4E96686B",
        521 => x"4E9CEBFF",
        522 => x"4EA36F08",
        523 => x"4EA9F188",
        524 => x"4EB0737E",
        525 => x"4EB6F4EA",
        526 => x"4EBD75CC",
        527 => x"4EC3F625",
        528 => x"4ECA75F5",
        529 => x"4ED0F53C",
        530 => x"4ED773F9",
        531 => x"4EDDF22D",
        532 => x"4EE46FD9",
        533 => x"4EEAECFC",
        534 => x"4EF16997",
        535 => x"4EF7E5A9",
        536 => x"4EFE6132",
        537 => x"4F04DC34",
        538 => x"4F0B56AE",
        539 => x"4F11D09F",
        540 => x"4F184A09",
        541 => x"4F1EC2EC",
        542 => x"4F253B46",
        543 => x"4F2BB31A",
        544 => x"4F322A66",
        545 => x"4F38A12B",
        546 => x"4F3F176A",
        547 => x"4F458D21",
        548 => x"4F4C0252",
        549 => x"4F5276FC",
        550 => x"4F58EB1F",
        551 => x"4F5F5EBC",
        552 => x"4F65D1D3",
        553 => x"4F6C4464",
        554 => x"4F72B66F",
        555 => x"4F7927F4",
        556 => x"4F7F98F4",
        557 => x"4F86096E",
        558 => x"4F8C7962",
        559 => x"4F92E8D2",
        560 => x"4F9957BB",
        561 => x"4F9FC620",
        562 => x"4FA63400",
        563 => x"4FACA15B",
        564 => x"4FB30E32",
        565 => x"4FB97A84",
        566 => x"4FBFE651",
        567 => x"4FC6519B",
        568 => x"4FCCBC5F",
        569 => x"4FD326A0",
        570 => x"4FD9905D",
        571 => x"4FDFF997",
        572 => x"4FE6624C",
        573 => x"4FECCA7E",
        574 => x"4FF3322C",
        575 => x"4FF99958",
        576 => x"50000000",
        577 => x"50066624",
        578 => x"500CCBC6",
        579 => x"501330E5",
        580 => x"50199582",
        581 => x"501FF99C",
        582 => x"50265D33",
        583 => x"502CC048",
        584 => x"503322DB",
        585 => x"503984EC",
        586 => x"503FE67A",
        587 => x"50464787",
        588 => x"504CA812",
        589 => x"5053081C",
        590 => x"505967A4",
        591 => x"505FC6AB",
        592 => x"50662530",
        593 => x"506C8334",
        594 => x"5072E0B8",
        595 => x"50793DBA",
        596 => x"507F9A3C",
        597 => x"5085F63D",
        598 => x"508C51BD",
        599 => x"5092ACBD",
        600 => x"5099073D",
        601 => x"509F613C",
        602 => x"50A5BABC",
        603 => x"50AC13BB",
        604 => x"50B26C3B",
        605 => x"50B8C43B",
        606 => x"50BF1BBC",
        607 => x"50C572BD",
        608 => x"50CBC93E",
        609 => x"50D21F41",
        610 => x"50D874C4",
        611 => x"50DEC9C8",
        612 => x"50E51E4E",
        613 => x"50EB7254",
        614 => x"50F1C5DC",
        615 => x"50F818E5",
        616 => x"50FE6B70",
        617 => x"5104BD7D",
        618 => x"510B0F0C",
        619 => x"5111601C",
        620 => x"5117B0AF",
        621 => x"511E00C3",
        622 => x"5124505A",
        623 => x"512A9F73",
        624 => x"5130EE0F",
        625 => x"51373C2D",
        626 => x"513D89CF",
        627 => x"5143D6F3",
        628 => x"514A2399",
        629 => x"51506FC3",
        630 => x"5156BB71",
        631 => x"515D06A1",
        632 => x"51635155",
        633 => x"51699B8C",
        634 => x"516FE547",
        635 => x"51762E86",
        636 => x"517C7749",
        637 => x"5182BF8F",
        638 => x"5189075A",
        639 => x"518F4EA9",
        640 => x"5195957C",
        641 => x"519BDBD3",
        642 => x"51A221AF",
        643 => x"51A86710",
        644 => x"51AEABF6",
        645 => x"51B4F060",
        646 => x"51BB344F",
        647 => x"51C177C4",
        648 => x"51C7BABD",
        649 => x"51CDFD3C",
        650 => x"51D43F41",
        651 => x"51DA80CA",
        652 => x"51E0C1DA",
        653 => x"51E7026F",
        654 => x"51ED428A",
        655 => x"51F3822B",
        656 => x"51F9C152",
        657 => x"52000000",
        658 => x"52063E33",
        659 => x"520C7BED",
        660 => x"5212B92D",
        661 => x"5218F5F5",
        662 => x"521F3242",
        663 => x"52256E17",
        664 => x"522BA972",
        665 => x"5231E455",
        666 => x"52381EBF",
        667 => x"523E58B0",
        668 => x"52449228",
        669 => x"524ACB28",
        670 => x"525103AF",
        671 => x"52573BBE",
        672 => x"525D7355",
        673 => x"5263AA74",
        674 => x"5269E11B",
        675 => x"5270174A",
        676 => x"52764D01",
        677 => x"527C8240",
        678 => x"5282B708",
        679 => x"5288EB59",
        680 => x"528F1F32",
        681 => x"52955293",
        682 => x"529B857E",
        683 => x"52A1B7F2",
        684 => x"52A7E9EE",
        685 => x"52AE1B74",
        686 => x"52B44C83",
        687 => x"52BA7D1C",
        688 => x"52C0AD3D",
        689 => x"52C6DCE9",
        690 => x"52CD0C1E",
        691 => x"52D33ADD",
        692 => x"52D96926",
        693 => x"52DF96F9",
        694 => x"52E5C456",
        695 => x"52EBF13D",
        696 => x"52F21DAE",
        697 => x"52F849AA",
        698 => x"52FE7530",
        699 => x"5304A041",
        700 => x"530ACADD",
        701 => x"5310F503",
        702 => x"53171EB5",
        703 => x"531D47F1",
        704 => x"532370B9",
        705 => x"5329990B",
        706 => x"532FC0E9",
        707 => x"5335E853",
        708 => x"533C0F48",
        709 => x"534235C8",
        710 => x"53485BD5",
        711 => x"534E816D",
        712 => x"5354A691",
        713 => x"535ACB41",
        714 => x"5360EF7D",
        715 => x"53671346",
        716 => x"536D369A",
        717 => x"5373597C",
        718 => x"53797BE9",
        719 => x"537F9DE4",
        720 => x"5385BF6B",
        721 => x"538BE07F",
        722 => x"5392011F",
        723 => x"5398214D",
        724 => x"539E4108",
        725 => x"53A46050",
        726 => x"53AA7F26",
        727 => x"53B09D89",
        728 => x"53B6BB79",
        729 => x"53BCD8F7",
        730 => x"53C2F603",
        731 => x"53C9129C",
        732 => x"53CF2EC4",
        733 => x"53D54A79",
        734 => x"53DB65BD",
        735 => x"53E1808F",
        736 => x"53E79AEF",
        737 => x"53EDB4DD",
        738 => x"53F3CE5A",
        739 => x"53F9E765",
        740 => x"54000000",
        741 => x"54061828",
        742 => x"540C2FE0",
        743 => x"54124727",
        744 => x"54185DFD",
        745 => x"541E7462",
        746 => x"54248A56",
        747 => x"542A9FDA",
        748 => x"5430B4ED",
        749 => x"5436C98F",
        750 => x"543CDDC1",
        751 => x"5442F183",
        752 => x"544904D5",
        753 => x"544F17B7",
        754 => x"54552A29",
        755 => x"545B3C2A",
        756 => x"54614DBC",
        757 => x"54675EDF",
        758 => x"546D6F91",
        759 => x"54737FD5",
        760 => x"54798FA8",
        761 => x"547F9F0D",
        762 => x"5485AE02",
        763 => x"548BBC88",
        764 => x"5491CA9F",
        765 => x"5497D847",
        766 => x"549DE581",
        767 => x"54A3F24B",
        768 => x"54A9FEA7",
        769 => x"54B00A94",
        770 => x"54B61613",
        771 => x"54BC2123",
        772 => x"54C22BC5",
        773 => x"54C835F9",
        774 => x"54CE3FBF",
        775 => x"54D44916",
        776 => x"54DA5200",
        777 => x"54E05A7C",
        778 => x"54E6628A",
        779 => x"54EC6A2A",
        780 => x"54F2715D",
        781 => x"54F87823",
        782 => x"54FE7E7B",
        783 => x"55048465",
        784 => x"550A89E3",
        785 => x"55108EF3",
        786 => x"55169397",
        787 => x"551C97CD",
        788 => x"55229B97",
        789 => x"55289EF3",
        790 => x"552EA1E4",
        791 => x"5534A467",
        792 => x"553AA67E",
        793 => x"5540A829",
        794 => x"5546A967",
        795 => x"554CAA39",
        796 => x"5552AA9F",
        797 => x"5558AA9A",
        798 => x"555EAA28",
        799 => x"5564A94A",
        800 => x"556AA800",
        801 => x"5570A64B",
        802 => x"5576A42A",
        803 => x"557CA19E",
        804 => x"55829EA6",
        805 => x"55889B43",
        806 => x"558E9774",
        807 => x"5594933B",
        808 => x"559A8E96",
        809 => x"55A08987",
        810 => x"55A6840C",
        811 => x"55AC7E27",
        812 => x"55B277D7",
        813 => x"55B8711C",
        814 => x"55BE69F7",
        815 => x"55C46268",
        816 => x"55CA5A6E",
        817 => x"55D05209",
        818 => x"55D6493B",
        819 => x"55DC4002",
        820 => x"55E23660",
        821 => x"55E82C53",
        822 => x"55EE21DD",
        823 => x"55F416FD",
        824 => x"55FA0BB3",
        825 => x"56000000",
        826 => x"5605F3E3",
        827 => x"560BE75C",
        828 => x"5611DA6D",
        829 => x"5617CD14",
        830 => x"561DBF52",
        831 => x"5623B126",
        832 => x"5629A292",
        833 => x"562F9395",
        834 => x"5635842F",
        835 => x"563B7460",
        836 => x"56416429",
        837 => x"56475389",
        838 => x"564D4281",
        839 => x"56533110",
        840 => x"56591F37",
        841 => x"565F0CF6",
        842 => x"5664FA4C",
        843 => x"566AE73B",
        844 => x"5670D3C1",
        845 => x"5676BFE0",
        846 => x"567CAB96",
        847 => x"568296E5",
        848 => x"568881CD",
        849 => x"568E6C4C",
        850 => x"56945665",
        851 => x"569A4016",
        852 => x"56A0295F",
        853 => x"56A61241",
        854 => x"56ABFABD",
        855 => x"56B1E2D1",
        856 => x"56B7CA7E",
        857 => x"56BDB1C4",
        858 => x"56C398A3",
        859 => x"56C97F1C",
        860 => x"56CF652E",
        861 => x"56D54AD9",
        862 => x"56DB301E",
        863 => x"56E114FD",
        864 => x"56E6F975",
        865 => x"56ECDD87",
        866 => x"56F2C132",
        867 => x"56F8A478",
        868 => x"56FE8758",
        869 => x"570469D1",
        870 => x"570A4BE5",
        871 => x"57102D93",
        872 => x"57160EDB",
        873 => x"571BEFBE",
        874 => x"5721D03B",
        875 => x"5727B053",
        876 => x"572D9005",
        877 => x"57336F53",
        878 => x"57394E3A",
        879 => x"573F2CBD",
        880 => x"57450ADB",
        881 => x"574AE894",
        882 => x"5750C5E8",
        883 => x"5756A2D7",
        884 => x"575C7F61",
        885 => x"57625B87",
        886 => x"57683748",
        887 => x"576E12A4",
        888 => x"5773ED9C",
        889 => x"5779C830",
        890 => x"577FA260",
        891 => x"57857C2B",
        892 => x"578B5593",
        893 => x"57912E96",
        894 => x"57970735",
        895 => x"579CDF71",
        896 => x"57A2B748",
        897 => x"57A88EBC",
        898 => x"57AE65CD",
        899 => x"57B43C79",
        900 => x"57BA12C3",
        901 => x"57BFE8A9",
        902 => x"57C5BE2B",
        903 => x"57CB934B",
        904 => x"57D16807",
        905 => x"57D73C60",
        906 => x"57DD1056",
        907 => x"57E2E3E9",
        908 => x"57E8B719",
        909 => x"57EE89E7",
        910 => x"57F45C52",
        911 => x"57FA2E5A",
        912 => x"58000000",
        913 => x"5805D143",
        914 => x"580BA223",
        915 => x"581172A2",
        916 => x"581742BE",
        917 => x"581D1278",
        918 => x"5822E1D0",
        919 => x"5828B0C6",
        920 => x"582E7F5A",
        921 => x"58344D8C",
        922 => x"583A1B5C",
        923 => x"583FE8CB",
        924 => x"5845B5D7",
        925 => x"584B8283",
        926 => x"58514ECD",
        927 => x"58571AB5",
        928 => x"585CE63C",
        929 => x"5862B162",
        930 => x"58687C27",
        931 => x"586E468A",
        932 => x"5874108D",
        933 => x"5879DA2E",
        934 => x"587FA36F",
        935 => x"58856C4E",
        936 => x"588B34CD",
        937 => x"5890FCEC",
        938 => x"5896C4AA",
        939 => x"589C8C07",
        940 => x"58A25304",
        941 => x"58A819A0",
        942 => x"58ADDFDC",
        943 => x"58B3A5B8",
        944 => x"58B96B34",
        945 => x"58BF304F",
        946 => x"58C4F50B",
        947 => x"58CAB967",
        948 => x"58D07D62",
        949 => x"58D640FE",
        950 => x"58DC043B",
        951 => x"58E1C717",
        952 => x"58E78994",
        953 => x"58ED4BB2",
        954 => x"58F30D70",
        955 => x"58F8CECF",
        956 => x"58FE8FCF",
        957 => x"5904506F",
        958 => x"590A10B0",
        959 => x"590FD092",
        960 => x"59159015",
        961 => x"591B4F39",
        962 => x"59210DFF",
        963 => x"5926CC65",
        964 => x"592C8A6D",
        965 => x"59324816",
        966 => x"59380561",
        967 => x"593DC24D",
        968 => x"59437EDB",
        969 => x"59493B0A",
        970 => x"594EF6DB",
        971 => x"5954B24E",
        972 => x"595A6D63",
        973 => x"59602819",
        974 => x"5965E272",
        975 => x"596B9C6D",
        976 => x"59715609",
        977 => x"59770F49",
        978 => x"597CC82A",
        979 => x"598280AE",
        980 => x"598838D4",
        981 => x"598DF09C",
        982 => x"5993A808",
        983 => x"59995F15",
        984 => x"599F15C6",
        985 => x"59A4CC19",
        986 => x"59AA820F",
        987 => x"59B037A8",
        988 => x"59B5ECE4",
        989 => x"59BBA1C3",
        990 => x"59C15646",
        991 => x"59C70A6B",
        992 => x"59CCBE34",
        993 => x"59D271A0",
        994 => x"59D824AF",
        995 => x"59DDD762",
        996 => x"59E389B8",
        997 => x"59E93BB2",
        998 => x"59EEED50",
        999 => x"59F49E91",
        1000 => x"59FA4F76",
        1001 => x"5A000000",
        1002 => x"5A05B02D",
        1003 => x"5A0B5FFE",
        1004 => x"5A110F73",
        1005 => x"5A16BE8C",
        1006 => x"5A1C6D49",
        1007 => x"5A221BAB",
        1008 => x"5A27C9B1",
        1009 => x"5A2D775C",
        1010 => x"5A3324AB",
        1011 => x"5A38D19E",
        1012 => x"5A3E7E36",
        1013 => x"5A442A73",
        1014 => x"5A49D655",
        1015 => x"5A4F81DB",
        1016 => x"5A552D07",
        1017 => x"5A5AD7D7",
        1018 => x"5A60824C",
        1019 => x"5A662C67",
        1020 => x"5A6BD626",
        1021 => x"5A717F8B",
        1022 => x"5A772895",
        1023 => x"5A7CD145"
    );
begin
    initial_guess_out <= INITIAL_GUESS_TABLE(to_integer(unsigned(address)));
end architecture;